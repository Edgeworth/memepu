`include "common.v"

module control_logic(
  input wire CLK,
  input wire N_CLK,
  input wire N_RST
);

  `ifdef FORMAL
  `endif
endmodule : control_logic
