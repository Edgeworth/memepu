`include "common.v"
module kpu(
  input wire CLK,
  input wire N_CLK,
  input wire N_RESET,
);

endmodule
